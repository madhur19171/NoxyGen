//`define VIVADO
//`define SHORTEST_PATH
`define XY
//`define VC
`define VC_DROP
//`define NO_VC
